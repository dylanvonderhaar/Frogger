module key_press_detector(

);


endmodule
